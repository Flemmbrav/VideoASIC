*****
***** Standards-compliant LVDS driver
*****
.SUBCKT LVDD D DGND VH Y0 Y1 VDD1 VSS
X1 DB N2  VDD1 DGND VSS inv4P
X2 D DB VDD1 DGND VSS inv4P
M1 N1 VH VDD1 VDD1 pch L=3u W=3.u M=100
M2 N1 N2 Y1 VSS nch L=0.4u W=1.2u M=40
M3 N1 DB Y0 VSS nch L=0.4u W=1.2u M=40
M4 Y1 DB CM VSS nch L=0.4u W=1.2u M=40
M5 Y0 N2 CM VSS nch L=0.4u W=1.2u M=40
M6 VDD1 VH VDD1 VDD1 pch L=3u W=3.u M=10
M7 CM CM DGND VSS nch  L=0.4u W=1.2u M=88
R7 Y1 Y0 10K TC=0.0, 0.0
.ENDS 
